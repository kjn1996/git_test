this is my code ....

version:0.02, this 's line is add in the version 0.02
