this is version 0.02 code txt
