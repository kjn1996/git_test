this is my code ....
